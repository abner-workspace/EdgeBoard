`timescale 1ns / 1ps
/****************************************************************
*   Auther : chengyang
*   Mail   : hn.cy@foxmail.com
*   Time   : 2019.09.06
*   Design :
*   Description :
*        PS write pL    ister
*    and PS read  PL    ister
*    Don't support busrt len, per transfer len = 1
****************************************************************/

module interconnect_stream
#(
    parameter  GP_ID_BITWIDTH                 = 4,
    parameter  GP_ADDR_BITWIDTH               = 32,
    parameter  GP_LEN_BITWIDTH                = 8,
    parameter  GP_SIZE_BITWIDTH               = 3,
    parameter  GP_BURST_BITWIDTH              = 2,
    parameter  GP_LOCK_BITWIDTH               = 1,
    parameter  GP_CACHE_BITWIDTH              = 4,
    parameter  GP_PROT_BITWIDTH               = 3,
    parameter  GP_QOS_BITWIDTH                = 4,
    parameter  GP_RESP_BITWIDTH               = 2,
    parameter  GP_DATA_BITWIDTH               = 32,
    parameter  GP_STRB_BITWIDTH               = GP_DATA_BITWIDTH/8,
    parameter  ARB_NUM                        = 1,
    parameter  PL_REGISTER_BASEADDR           = 32'h0000_0000,
    parameter  PS_REGISTER_BASEADDR           = 32'h0000_0000
)(
    input                                       sys_clk,
    input                                       sys_rst,
// config PL
    input       [GP_ID_BITWIDTH-1 : 0]          s_axi_awid,
    input       [GP_ADDR_BITWIDTH-1 : 0]        s_axi_awaddr,
    input       [GP_LEN_BITWIDTH-1 : 0]         s_axi_awlen,
    input       [GP_SIZE_BITWIDTH-1 : 0]        s_axi_awsize,
    input       [GP_BURST_BITWIDTH-1 : 0]       s_axi_awburst,
    input       [GP_LOCK_BITWIDTH-1 : 0]        s_axi_awlock,
    input       [GP_CACHE_BITWIDTH-1 : 0]       s_axi_awcache,
    input       [GP_PROT_BITWIDTH-1 : 0]        s_axi_awprot,
    input       [GP_QOS_BITWIDTH-1 : 0]         s_axi_awqos,
    input                                       s_axi_awvalid,
    output                                      s_axi_awready,
    input       [GP_ID_BITWIDTH-1 : 0]          s_axi_wid,
    input       [GP_DATA_BITWIDTH-1 : 0]        s_axi_wdata,
    input       [GP_STRB_BITWIDTH-1 : 0]        s_axi_wstrb,
    input                                       s_axi_wlast,
    input                                       s_axi_wvalid,
    output                                      s_axi_wready,
    output      [GP_ID_BITWIDTH-1 : 0]          s_axi_bid,
    output      [GP_RESP_BITWIDTH-1 : 0]        s_axi_bresp,
    output                                      s_axi_bvalid,
    input                                       s_axi_bready,
    input       [GP_PROT_BITWIDTH-1 : 0]        s_axi_arprot,
    input       [GP_ID_BITWIDTH-1 : 0]          s_axi_arid,
    input       [GP_ADDR_BITWIDTH-1 : 0]        s_axi_araddr,
    input       [GP_LEN_BITWIDTH-1 : 0]         s_axi_arlen,
    input       [GP_SIZE_BITWIDTH-1 : 0]        s_axi_arsize,
    input       [GP_BURST_BITWIDTH-1 : 0]       s_axi_arburst,
    input       [GP_LOCK_BITWIDTH-1 : 0]        s_axi_arlock,
    input       [GP_CACHE_BITWIDTH-1 : 0]       s_axi_arcache,
    input       [GP_QOS_BITWIDTH-1 : 0]         s_axi_arqos,
    input                                       s_axi_arvalid,
    output                                      s_axi_arready,
    output      [GP_ID_BITWIDTH-1 : 0]          s_axi_rid,
    output      [GP_DATA_BITWIDTH-1 : 0]        s_axi_rdata,
    output      [GP_RESP_BITWIDTH-1 : 0]        s_axi_rresp,
    output                                      s_axi_rlast,
    output                                      s_axi_rvalid,
    input                                       s_axi_rready,
// config PS
    output      [GP_ID_BITWIDTH-1 : 0]          m_axi_awid,
    output      [GP_ADDR_BITWIDTH-1 : 0]        m_axi_awaddr,
    output      [GP_LEN_BITWIDTH-1 : 0]         m_axi_awlen,
    output      [GP_SIZE_BITWIDTH-1 : 0]        m_axi_awsize,
    output      [GP_BURST_BITWIDTH-1 : 0]       m_axi_awburst,
    output      [GP_LOCK_BITWIDTH-1 : 0]        m_axi_awlock,
    output      [GP_CACHE_BITWIDTH-1 : 0]       m_axi_awcache,
    output      [GP_PROT_BITWIDTH-1 : 0]        m_axi_awprot,
    output      [GP_QOS_BITWIDTH-1 : 0]         m_axi_awqos,
    output                                      m_axi_awvalid,
    input                                       m_axi_awready,
    output      [GP_ID_BITWIDTH-1 : 0]          m_axi_wid,
    output      [GP_DATA_BITWIDTH-1 : 0]        m_axi_wdata,
    output      [GP_STRB_BITWIDTH-1 : 0]        m_axi_wstrb,
    output                                      m_axi_wlast,
    output                                      m_axi_wvalid,
    input                                       m_axi_wready,
    input       [GP_ID_BITWIDTH-1 : 0]          m_axi_bid,
    input       [GP_RESP_BITWIDTH-1 : 0]        m_axi_bresp,
    input                                       m_axi_bvalid,
    output                                      m_axi_bready,
    output      [GP_PROT_BITWIDTH-1 : 0]        m_axi_arprot,
    output      [GP_ID_BITWIDTH-1 : 0]          m_axi_arid,
    output      [GP_ADDR_BITWIDTH-1 : 0]        m_axi_araddr,
    output      [GP_LEN_BITWIDTH-1 : 0]         m_axi_arlen,
    output      [GP_SIZE_BITWIDTH-1 : 0]        m_axi_arsize,
    output      [GP_BURST_BITWIDTH-1 : 0]       m_axi_arburst,
    output      [GP_LOCK_BITWIDTH-1 : 0]        m_axi_arlock,
    output      [GP_CACHE_BITWIDTH-1 : 0]       m_axi_arcache,
    output      [GP_QOS_BITWIDTH-1 : 0]         m_axi_arqos,
    output                                      m_axi_arvalid,
    input                                       m_axi_arready,
    input       [GP_ID_BITWIDTH-1 : 0]          m_axi_rid,
    input       [GP_DATA_BITWIDTH-1 : 0]        m_axi_rdata,
    input       [GP_RESP_BITWIDTH-1 : 0]        m_axi_rresp,
    input                                       m_axi_rlast,
    input                                       m_axi_rvalid,
    output                                      m_axi_rready,
// register
    output                                      upload_result_next,
    input                                       upload_result_en,
    input       [31 : 0]                        upload_result_addr,
    input       [31 : 0]                        upload_result_nbyte,
    output      [31 : 0]                        update_status,
    input       [31 : 0]                        set_arg_std,
    output                                      platform_init_done,
    output      [7 : 0]                         sdi_sync_std,
    input       [31 : 0]                        sys_uhdsdi_status,
    output                                      sys_uhdsdi_soft_rst,
    output                                      sys_hdmi_soft_rst,
    output      [31 : 0]                        sys_device_id1,
    output      [31 : 0]                        sys_device_id2,
    output      [31 : 0]                        sys_device_id3,
    output      [31 : 0]                        sys_device_id4,
    output      [31 : 0]                        sys_device_arg1,
    input       [12*8-1 : 0]                    sys_device_mac,
// user define interface
    // write
    output  [ARB_NUM*1-1 : 0]                   write_cmd_done,
    input   [ARB_NUM*1-1 : 0]                   write_cmd_start,
    input   [ARB_NUM*GP_ADDR_BITWIDTH-1 : 0]    write_cmd_addr,
    input   [ARB_NUM*GP_ADDR_BITWIDTH-1 : 0]    write_cmd_len,
    output  [ARB_NUM*1-1 : 0]                   write_axis_ready,
    input   [ARB_NUM*1-1 : 0]                   write_axis_valid,
    input   [ARB_NUM*GP_DATA_BITWIDTH-1 : 0]    write_axis_data,
    input   [ARB_NUM*GP_STRB_BITWIDTH-1 : 0]    write_axis_strb,
    input   [ARB_NUM*1-1 : 0]                   write_axis_last,
    // read
    output  [ARB_NUM*1-1 : 0]                   read_cmd_done,
    input   [ARB_NUM*1-1 : 0]                   read_cmd_start,
    input   [ARB_NUM*GP_ADDR_BITWIDTH-1 : 0]    read_cmd_addr,
    input   [ARB_NUM*GP_ADDR_BITWIDTH-1 : 0]    read_cmd_len,
    input   [ARB_NUM*1-1 : 0]                   read_axis_ready,
    output  [ARB_NUM*1-1 : 0]                   read_axis_valid,
    output  [ARB_NUM*GP_DATA_BITWIDTH-1 : 0]    read_axis_data,
    output  [ARB_NUM*1-1 : 0]                   read_axis_last
);


config_pl_register #(
    .GP_ID_BITWIDTH                 (GP_ID_BITWIDTH),
    .GP_ADDR_BITWIDTH               (GP_ADDR_BITWIDTH),
    .GP_LEN_BITWIDTH                (GP_LEN_BITWIDTH),
    .GP_SIZE_BITWIDTH               (GP_SIZE_BITWIDTH),
    .GP_BURST_BITWIDTH              (GP_BURST_BITWIDTH),
    .GP_LOCK_BITWIDTH               (GP_LOCK_BITWIDTH),
    .GP_CACHE_BITWIDTH              (GP_CACHE_BITWIDTH),
    .GP_PROT_BITWIDTH               (GP_PROT_BITWIDTH),
    .GP_QOS_BITWIDTH                (GP_QOS_BITWIDTH),
    .GP_RESP_BITWIDTH               (GP_RESP_BITWIDTH),
    .GP_DATA_BITWIDTH               (GP_DATA_BITWIDTH),
    .GP_STRB_BITWIDTH               (GP_STRB_BITWIDTH),
    .REGISTER_BASEADDR              (PL_REGISTER_BASEADDR)
) inst_config_pl_register (
    .sys_clk                        (sys_clk),
    .sys_rst                        (sys_rst),
    .s_axi_awid                     (s_axi_awid),
    .s_axi_awaddr                   (s_axi_awaddr),
    .s_axi_awlen                    (s_axi_awlen),
    .s_axi_awsize                   (s_axi_awsize),
    .s_axi_awburst                  (s_axi_awburst),
    .s_axi_awlock                   (s_axi_awlock),
    .s_axi_awcache                  (s_axi_awcache),
    .s_axi_awprot                   (s_axi_awprot),
    .s_axi_awqos                    (s_axi_awqos),
    .s_axi_awvalid                  (s_axi_awvalid),
    .s_axi_awready                  (s_axi_awready),
    .s_axi_wid                      (s_axi_wid),
    .s_axi_wdata                    (s_axi_wdata),
    .s_axi_wstrb                    (s_axi_wstrb),
    .s_axi_wlast                    (s_axi_wlast),
    .s_axi_wvalid                   (s_axi_wvalid),
    .s_axi_wready                   (s_axi_wready),
    .s_axi_bid                      (s_axi_bid),
    .s_axi_bresp                    (s_axi_bresp),
    .s_axi_bvalid                   (s_axi_bvalid),
    .s_axi_bready                   (s_axi_bready),
    .s_axi_arprot                   (s_axi_arprot),
    .s_axi_arid                     (s_axi_arid),
    .s_axi_araddr                   (s_axi_araddr),
    .s_axi_arlen                    (s_axi_arlen),
    .s_axi_arsize                   (s_axi_arsize),
    .s_axi_arburst                  (s_axi_arburst),
    .s_axi_arlock                   (s_axi_arlock),
    .s_axi_arcache                  (s_axi_arcache),
    .s_axi_arqos                    (s_axi_arqos),
    .s_axi_arvalid                  (s_axi_arvalid),
    .s_axi_arready                  (s_axi_arready),
    .s_axi_rid                      (s_axi_rid),
    .s_axi_rdata                    (s_axi_rdata),
    .s_axi_rresp                    (s_axi_rresp),
    .s_axi_rlast                    (s_axi_rlast),
    .s_axi_rvalid                   (s_axi_rvalid),
    .s_axi_rready                   (s_axi_rready),
// PL Register
    .upload_result_next             (upload_result_next),
    .upload_result_en               (upload_result_en),
    .upload_result_addr             (upload_result_addr),
    .upload_result_nbyte            (upload_result_nbyte),
    .update_status                  (update_status),
    .set_arg_std                    (set_arg_std),
    .platform_init_done             (platform_init_done),
    .sdi_sync_std                   (sdi_sync_std),
    .sys_uhdsdi_status              (sys_uhdsdi_status),
    .sys_uhdsdi_soft_rst            (sys_uhdsdi_soft_rst),
    .sys_hdmi_soft_rst              (sys_hdmi_soft_rst),
    .sys_device_id1                 (sys_device_id1),
    .sys_device_id2                 (sys_device_id2),
    .sys_device_id3                 (sys_device_id3),
    .sys_device_id4                 (sys_device_id4),
    .sys_device_arg1                (sys_device_arg1),
    .sys_device_mac                 (sys_device_mac)
);

axi_arb_interface #(
    .AXI_ID_BITWIDTH        (GP_ID_BITWIDTH),
    .AXI_ADDR_BITWIDTH      (GP_ADDR_BITWIDTH),
    .AXI_LEN_BITWIDTH       (GP_LEN_BITWIDTH),
    .AXI_SIZE_BITWIDTH      (GP_SIZE_BITWIDTH),
    .AXI_BURST_BITWIDTH     (GP_BURST_BITWIDTH),
    .AXI_LOCK_BITWIDTH      (GP_LOCK_BITWIDTH),
    .AXI_CACHE_BITWIDTH     (GP_CACHE_BITWIDTH),
    .AXI_PROT_BITWIDTH      (GP_PROT_BITWIDTH),
    .AXI_QOS_BITWIDTH       (GP_QOS_BITWIDTH),
    .AXI_RESP_BITWIDTH      (GP_RESP_BITWIDTH),
    .AXI_DATA_BITWIDTH      (GP_DATA_BITWIDTH),
    .AXI_STRB_BITWIDTH      (GP_STRB_BITWIDTH),
    .BURST_MAX              (16),
    .ARB_NUM                (1),
    .ID                     (0)
) inst_config_ps_register (
    .sys_clk                (sys_clk),
    .sys_rst                (sys_rst),
    .write_cmd_done         (write_cmd_done),
    .write_cmd_start        (write_cmd_start),
    .write_cmd_addr         (write_cmd_addr),
    .write_cmd_len          (write_cmd_len),
    .write_axis_ready       (write_axis_ready),
    .write_axis_valid       (write_axis_valid),
    .write_axis_data        (write_axis_data),
    .write_axis_strb        (8'hFF),
    .write_axis_last        (write_axis_last),
    .read_cmd_done          (),
    .read_cmd_start         (0),
    .read_cmd_addr          (),
    .read_cmd_len           (),
    .read_axis_ready        (),
    .read_axis_valid        (),
    .read_axis_data         (),
    .read_axis_last         (),
    .m_axi_awid             (m_axi_awid),
    .m_axi_awaddr           (m_axi_awaddr),
    .m_axi_awlen            (m_axi_awlen),
    .m_axi_awsize           (m_axi_awsize),
    .m_axi_awburst          (m_axi_awburst),
    .m_axi_awlock           (m_axi_awlock),
    .m_axi_awcache          (m_axi_awcache),
    .m_axi_awprot           (m_axi_awprot),
    .m_axi_awqos            (m_axi_awqos),
    .m_axi_awvalid          (m_axi_awvalid),
    .m_axi_awready          (m_axi_awready),
    .m_axi_wid              (m_axi_wid),
    .m_axi_wdata            (m_axi_wdata),
    .m_axi_wstrb            (m_axi_wstrb),
    .m_axi_wlast            (m_axi_wlast),
    .m_axi_wvalid           (m_axi_wvalid),
    .m_axi_wready           (m_axi_wready),
    .m_axi_bid              (m_axi_bid),
    .m_axi_bresp            (m_axi_bresp),
    .m_axi_bvalid           (m_axi_bvalid),
    .m_axi_bready           (m_axi_bready),
    .m_axi_arid             (m_axi_arid),
    .m_axi_araddr           (m_axi_araddr),
    .m_axi_arlen            (m_axi_arlen),
    .m_axi_arsize           (m_axi_arsize),
    .m_axi_arburst          (m_axi_arburst),
    .m_axi_arlock           (m_axi_arlock),
    .m_axi_arcache          (m_axi_arcache),
    .m_axi_arprot           (m_axi_arprot),
    .m_axi_arqos            (m_axi_arqos),
    .m_axi_arvalid          (m_axi_arvalid),
    .m_axi_arready          (m_axi_arready),
    .m_axi_rid              (m_axi_rid),
    .m_axi_rdata            (m_axi_rdata),
    .m_axi_rresp            (m_axi_rresp),
    .m_axi_rlast            (m_axi_rlast),
    .m_axi_rvalid           (m_axi_rvalid),
    .m_axi_rready           (m_axi_rready)
);

endmodule